library verilog;
use verilog.vl_types.all;
entity FSM_vlg_check_tst is
    port(
        done            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FSM_vlg_check_tst;
